module (
    input button1,
    input button2
)
endmodle

///new